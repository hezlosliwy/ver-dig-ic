package vdic_dut_2023_pkg;
	
import misc_pkg::*;
`include "coverage.svh"
`include "tpgen.svh"
`include "scoreboard.svh"
`include "testbench.svh"

endpackage