//----------------------------------------------------------------------
// Created by Stanislaw Klat on Wed Jan 03 20:41:39 CET 2024
//----------------------------------------------------------------------

//This is a dummy DUT.
module dut(
    input wire clock,
    input wire reset,
    input wire [32:0] data
  );

endmodule : dut
