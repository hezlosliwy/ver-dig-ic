package vdic_dut_2023_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import misc_pkg::*;
`include "random_command.svh"
`include "minmax_command.svh"
`include "result_transaction.svh"
`include "coverage.svh"
`include "scoreboard.svh"
`include "driver.svh"
`include "data_monitor.svh"
`include "result_monitor.svh"
`include "tpgen.svh"
`include "env.svh"
`include "random_test.svh"
`include "min_max_test.svh"


endpackage