package vdic_dut_2023_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import misc_pkg::*;
`include "vdic_dut_2023_agent_config.svh"
`include "random_command.svh"
`include "minmax_command.svh"
`include "stim_module.svh"
`include "result_transaction.svh"
`include "coverage.svh"
`include "scoreboard.svh"
`include "driver.svh"
`include "data_monitor.svh"
`include "result_monitor.svh"
`include "tpgen.svh"

`include "vdic_dut_2023_agent.svh"

`include "env_config.svh"
`include "env.svh"
`include "dual_test.svh"

endpackage