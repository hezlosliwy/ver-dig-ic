package shapes_pkg;
	`include "shape_c.svh"
	`include "circle_c.svh"
	`include "rectangle_c.svh"
	`include "triangle_c.svh"
	`include "polygon_c.svh"
endpackage