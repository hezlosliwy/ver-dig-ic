package vdic_dut_2023_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import misc_pkg::*;
`include "coverage.svh"
`include "scoreboard.svh"
`include "driver.svh"
`include "data_monitor.svh"
`include "result_monitor.svh"
`include "base_tpgen.svh"
`include "random_tpgen.svh"
`include "min_max_tpgen.svh"
`include "env.svh"
`include "random_test.svh"
`include "min_max_test.svh"


endpackage