package shape_pkg;

    typedef struct {
        real x;
        real y;
    } point;

	typedef enum {CIRCLE, TRIANGLE, RECTANGLE, POLYGON, NO_SHAPE} e_shape;

endpackage