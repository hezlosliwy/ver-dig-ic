//----------------------------------------------------------------------
// Created by Stanislaw Klat on Wed Jan 03 20:41:39 CET 2024
//----------------------------------------------------------------------

package sk_test_pkg;

  `include "uvm_macros.svh"
  import uvm_pkg::*;

  import sk_pkg::*;

  // HINT Here you include tests.

  `include "sk_base_test.svh"
  `include "sk_example_test.svh"


endpackage : sk_test_pkg
