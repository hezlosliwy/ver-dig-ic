package shape_pkg;

    typedef struct {
        real x;
        real y;
    } point;

endpackage